module FSMPaceMaker ();

endmodule

