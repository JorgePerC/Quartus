// #Import MUX, PROCESSOR REGISTER
// No need to import, since all the files were overwitten

module CPU ();


endmodule
