
`timescale 1ns / 1ps


module Mux8_test;

	reg [7:0] A;
	reg [7:0] B;
	reg [7:0] C;
	reg [7:0] D;
	reg [7:0] E;
	reg [7:0] F;
	reg [7:0] G;
	reg [7:0] H;
	reg [2:0] S; // 2 pq log2(8) = 3 | 3-1 0 2

	wire [7:0] OUT;

	Mux8 uut (
		.A(A),
		.B(B),
		.C(C),
		.D(D),
		.E(E),
		.F(F),
		.G(G),
		.H(H),
		.S(S),
		.OUT (OUT)
	
	);

initial begin 

// 1
A = 0;
	B = 0;
	C = 0;
	D = 1;
	E = 0;
	F = 0;
	G = 0;
	H = 0;
	S = 0;

	#10;

// 2
A = 9;
	B = 10;
	C = 131;
	D = 15;
	E = 150;
	F = 21;
	G = 50;
	H = 200;
	S = 1;

	#10;

//3
A = 9;
	B = 103;
	C = 101;
	D = 157;
	E = 150;
	F = 20;
	G = 50;
	H = 200;
	S = 2;

	#10;

//4
A = 9;
	B = 17;
	C = 101;
	D = 15;
	E = 150;
	F = 20;
	G = 60;
	H = 200;
	S = 3;

	#10;

//5
A = 99;
	B = 10;
	C = 101;
	D = 15;
	E = 150;
	F = 20;
	G = 50;
	H = 200;
	S = 4;

	#10;
//6
A = 95;
	B = 10;
	C = 101;
	D = 15;
	E = 180;
	F = 20;
	G = 50;
	H = 200;
	S = 5;
	
	#10;
//7
A = 91;
	B = 10;
	C = 101;
	D = 15;
	E = 150;
	F = 20;
	G = 50;
	H = 210;
	S = 6;
	#10;

//8
A = 19;
	B = 10;
	C = 11;
	D = 15;
	E = 150;
	F = 20;
	G = 57;
	H = 200;
	S = 7;

	#10;

//9
A = 59;
	B = 20;
	C = 101;
	D = 154;
	E = 150;
	F = 20;
	G = 57;
	H = 200;
	S = 7;
	#10;
// 10
A = 30;
	B = 0;
	C = 6;
	D = 23;
	E = 54;
	F = 58;
	G = 78;
	H = 107;
	S = 150;

	#10;
// 11
A = 50;
	B = 0;
	C = 0;
	D = 0;
	E = 0;
	F = 0;
	G = 0;
	H = 0;
	S = 0;

	#10;

// 12
A = 7;
	B = 50;
	C = 101;
	D = 35;
	E = 150;
	F = 20;
	G = 50;
	H = 200;
	S = 1;

	#10;

//13
A = 9;
	B = 10;
	C = 41;
	D = 155;
	E = 150;
	F = 20;
	G = 150;
	H = 200;
	S = 23;

	#10;

//14
A = 9;
	B = 15;
	C = 101;
	D = 75;
	E = 150;
	F = 27;
	G = 50;
	H = 200;
	S = 3;

	#10;

//15
A = 8;
	B = 10;
	C = 11;
	D = 65;
	E = 150;
	F = 80;
	G = 59;
	H = 200;
	S = 4;

	#10;

//16
A = 35;
	B = 106;
	C = 121;
	D = 13;
	E = 150;
	F = 27;
	G = 50;
	H = 200;
	S = 5;
	#10;
//17
A = 9;
	B = 10;
	C = 101;
	D = 157;
	E = 10;
	F = 2;
	G = 57;
	H = 20;
	S = 65;
	#10;
//18
A = 92;
	B = 40;
	C = 101;
	D = 13;
	E = 150;
	F = 27;
	G = 50;
	H = 200;
	S = 7;
	#10;
//19
A = 9;
	B = 10;
	C = 101;
	D = 15;
	E = 150;
	F = 20;
	G = 50;
	H = 200;
	S = 7;
	#10;
// 20
A = 5;
	B = 0;
	C = 34;
	D = 0;
	E = 0;
	F = 45;
	G = 0;
	H = 0;
	S = 7;

	#10;
// 21
A = 50;
	B = 34;
	C = 0;
	D = 5;
	E = 23;
	F = 0;
	G = 67;
	H = 0;
	S = 0;

	#10;

// 22
A = 9;
	B = 10;
	C = 101;
	D = 15;
	E = 150;
	F = 20;
	G = 50;
	H = 200;
	S = 1;

	#10;

//23
A = 57;
	B = 16;
	C = 161;
	D = 15;
	E = 150;
	F = 23;
	G = 50;
	H = 200;
	S = 2;

	#10;

//24
A = 45;
	B = 10;
	C = 141;
	D = 5;
	E = 150;
	F = 20;
	G = 53;
	H = 200;
	S = 3;

	#10;

end
endmodule

