module PaceMakerCool (

);
// Timer (contador) 
// FSM


endmodule