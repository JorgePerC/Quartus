//Import processor register 

module MemoryRegister ();

endmodule
