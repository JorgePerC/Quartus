// TODO: DELETE THIS.
module ALU ();

endmodule
