module FSMPaceMaker ();

endmodule
