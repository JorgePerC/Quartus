module PaceMaker (

);
// Timer (contador) 
// FSM


endmodule
